/*
 * Current working ALU design for Group 9 
 * Group Members: Ben Leaptrot, Christian Giauque, Colton Watson, Nathan Hummel
 *
 * Last updated: September 7, 2020
 *
 * Inputs: 
 *   A: Source A - 16-bit value
 *   B: Source B - 16-bit value
 *   Opcode: 8-bit opcode designating which instruction to execute
 *
 * Outputs:
 *   C: 16-bit value from opcode computation.
 *   Flags: 5-bit array of bits. 1=true, 0=false. The bits currently correspond to these flags:
 *            Carry flag    (carry/borrow from addition/subtraction) - Bit 4
 *            Low flag      (unsigned integer comparison)            - Bit 3
 *            Overflow flag (signed arithmetic overflow)             - Bit 2
 *            Zero flag     (operation left zero in the output)      - Bit 1
 *            Negative flag (signed integer comparison)              - Bit 0
 *
 * Notes:
 *   Baseline Operations not currently implemented (I'm not sure how yet): LOAD, STOR, BCOND, JCOND, JAL
 *   Is the borrow flag correctly set in the subtraction operations?
 *   Are logical/arithmetic shifts incorporated correctly?
 *     arithmetic shifts aren't baseline, but are highly recommneded (commented out right now)
 * 
 */
module alu(A, B, C, Opcode, Flags);

	input  [15:0] A, B;
	input  [7:0]  Opcode;
	
	output reg [15:0] C;
	output reg [4:0]  Flags;
	
	// Flags
	parameter carry_f    = 3'd4;
	parameter low_f      = 3'd3;
	parameter overflow_f = 3'd2;
	parameter zero_f     = 3'd1;
	parameter negative_f = 3'd0;

	// Opcodes
	// * = Baseline instructions
	// Obviously delete unused/unneeded parameters.
	parameter ADD  = 8'b00000101; // *
	parameter ADDI = 8'b0101xxxx; // *
	parameter ADDU = 8'b00000110;
	parameter ADDUI= 8'b0110xxxx;
	parameter ADDC = 8'b00000111;
	parameter ADDCI= 8'b0111xxxx;
	
	parameter SUB  = 8'b00001001; // *
	parameter SUBI = 8'b1001xxxx; // *
	parameter SUBC = 8'b00001010;
	parameter SUBCI= 8'b1010xxxx; 
	parameter CMP  = 8'b00001011; // *
	parameter CMPI = 8'b1011xxxx; // *
	parameter AND  = 8'b00000001; // *
	parameter ANDI = 8'b0001xxxx; // *
	parameter OR   = 8'b00000010; // *
	parameter ORI  = 8'b0010xxxx; // *
	parameter XOR  = 8'b00000011; // *
	parameter XORI = 8'b0011xxxx; // *
	parameter MOV  = 8'b00001101; // *
	parameter MOVI = 8'b1101xxxx; // *
	parameter LSH  = 8'b10000100; // *
	parameter LSHI = 8'b1000000x; // x -> sign (0=left, 2's comp)
	parameter ASHU = 8'b10000110;
	parameter ASHUI= 8'b1000001x; // x -> sign (0=left, 2's comp)
	parameter LUI  = 8'b1111xxxx; // *
	
	/* How should these be done in the ALU? */
	parameter LOAD = 8'b01000000; // *
	parameter STOR = 8'b01000100; // *
	parameter Bcond= 8'b1100xxxx; // *
	parameter Jcond= 8'b01001100; // *
	parameter JAL  = 8'b01001000; // *
	
	
	always@(A, B, Opcode)
	begin		
		
		Flags = 5'b0;
		C = 16'b0;
		
		casex (Opcode)
		ADD: // Integer addition
			begin
			{Flags[carry_f], C} = A + B; 
			
			// Overflow occurs when (pos) + (pos) = neg
			//             and when (neg) + (neg) = pos
			if((~A[15] & ~B[15] & C[15]) | (A[15] & B[15] & ~C[15])) 
				Flags[overflow_f] = 1'b1;
			end
			
		ADDI: // Integer addition immediate
			begin
			// B is thought of as being an 8-bit number, sign-extend it.
			{Flags[carry_f], C} = A + {{8{B[7]}} , B[7:0]};
			
			if((~A[15] & ~B[15] & C[15]) | (A[15] & B[15] & ~C[15])) 
				Flags[overflow_f] = 1'b1;
			end
			
		ADDU: // Integer addition, no flags will be set
			begin
			C = A + B; 
			end
			
		SUB: // Integer subtraction
			begin
			{Flags[carry_f], C} = A - B;
			
			if(A == B) 
				Flags[zero_f] = 1'b1; 
			
			// Overflow occurs when (pos) - (neg) = neg
			//             and when (neg) - (pos) = pos
			if((A[15] & ~B[15] & ~C[15]) | (~A[15] & B[15] & C[15])) 
				Flags[overflow_f] = 1'b1;
			
			if(A < B)
				Flags[low_f] = 1'b1;
				
			if($signed(A) < $signed(B))
				Flags[negative_f] = 1'b1;			
			
			end
			
		SUBI: // Integer subtraction immediate
			begin
			{Flags[carry_f], C} = A - {{8{B[7]}} , B[7:0]};
			
			if(A == B) 
				Flags[zero_f] = 1'b1; 
			
			if((A[15] & ~B[7] & ~C[15]) | (~A[15] & B[7] & C[15])) 
				Flags[overflow_f] = 1'b1;
			
			if(A < B)
				Flags[low_f] = 1'b1;
			
			if($signed(A) < $signed(B))
				Flags[negative_f] = 1'b1;
			
			end
		
		CMP: // Comparison. Affects PSR.Z, PSR.N, PSR.L.
			begin
			
			if(A == B)
				Flags[zero_f] = 1'b1;
				
			if($signed(A) < $signed(B))
				Flags[negative_f] = 1'b1;
				
			if(A < B)
				Flags[low_f] = 1'b1;
			
			end
			
		CMPI: // Comparison immediate
			begin 
			if(A == {{8{B[7]}} , B[7:0]})
				Flags[zero_f] = 1'b1;
				
			if($signed(A) < $signed({{8{B[7]}} , B[7:0]}))
				Flags[negative_f] = 1'b1;
				
			if(A < {8'b0 , B[7:0]})
				Flags[low_f] = 1'b1;
			end

		AND: // Logical AND
			begin
			C = A & B;
			
			if(C == 16'b0)
				Flags[zero_f] = 1'b1;
			end
			
		ANDI: // Logical AND with zero-extended immediate
			begin
			C = A & {8'b0 , B[7:0]}; 
			
			if(C == 16'b0)
				Flags[zero_f] = 1'b1;
			end
			
		OR: // Logical OR
			begin
			C = A | B; 
			end
			
		ORI: // Logical OR with zero-extended immediate
			begin
			C = A | {8'b0 , B[7:0]}; 
			end
			
		XOR: // Logical XOR 
			begin
			C = A ^ B;
			end
			
		XORI: // Logical XOR with zero-extended immediate
			begin
			C = A ^ {8'b0 , B[7:0]}; 
			end
			
		MOV: // Move
			begin
			C = B; 
			end
			
		MOVI: // Move with zero-extended immediate 
			begin
			C = {8'b0 , B[7:0]}; 
			end
			
		LSH: // Logical Shift
			begin
			C = A << B; // Need to check if B is weird?
			end
			
		LSHI:
			begin
			if(Opcode[0] == 1'b0)
				begin
				C = A << B;
				//C = A << $signed(B[5:0]); // <- Do it like that?
				end
			else
				begin
				C = A <<< B;
				end
			end
			/*
		ASHU: // Arithmetic Shift
			begin
			C = A <<< B;
			end
		ASHUI:
			begin
			C = A <<< B;
			end
			*/
		LUI: // Load upper immediate (Move, but fill MSB with immediate)
			begin
			C = {B [7:0], 8'b0}; 
			end
//		LOAD: // Load from Memory
//			begin
//			C = mem[B]; // ???
//			end
//    STOR: // Store in memory
//			begin
//			// mem[A] = B; ???
//			end
//		Bcond:
//			begin
//       // A = COND
//       // 
//			PC - $signed(
//			end
//		Jcond:
//			begin
//			end
//		JAL:
//			begin
//			end
		
		default:
			begin
				C = 16'b0;
				Flags = 5'b0;
			end		
		endcase
		
	end
	
endmodule
