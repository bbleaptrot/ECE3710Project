module fsm(clk, rst, PCen, Ren, RegOrImm);
input clk, rst;
output PCen, RegOrImm;
output [15:0] Ren;

endmodule